//Jorge Avila Juarez 1001543128
module CLA (
inout AddSub,
input [7:0] A,B,
output [7:0] R,
output Cout,
output OVR);



endmodule 