module KnightRiderFlasher(





);

endmodule
